package router_pkg;
import uvm_pkg::*;
`include "uvm_macros.svh"

`include "source_xtn.sv"
`include "corrupt_source_xtn.sv"

`include "dest_xtn.sv"
`include "source_config.sv"
`include "dest_config.sv"
`include "tb_config.sv"

`include "source_driver.sv"
`include "source_monitor.sv"
`include "source_sequencer.sv"

`include "dest_driver.sv"
`include "dest_sequencer.sv"
`include "dest_monitor.sv"

`include "source_agent.sv"
`include "dest_agent.sv"

`include "source_agent_top.sv"
`include "dest_agent_top.sv"
`include "virtual_sequencer.sv"

`include "router_sb.sv"
`include "env.sv"

`include "source_seqs.sv"
`include "dest_seqs.sv"

`include "virtual_sequence.sv"
`include "test.sv"

endpackage
